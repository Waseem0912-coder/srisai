skdfjlksdfjskadfj:

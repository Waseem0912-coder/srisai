skdfjlksdfjskadfj:
werwker
